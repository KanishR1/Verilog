module xor_gate (
    input A,B, output S
);
assign S = A^B;
    
endmodule